--Component.vhdl
--設計名稱 | Design name
--	
--更新紀錄 | Changelog
--	Changelog is now stored on GitHub(http://www.github.com)
--已知問題 | Known issues
--	Known issues is now stored on GitHub(http://www.github.com)
--待辦事項 | Todos
--	Todo is now stored on GitHub(http://www.github.com)
--著作權宣告 | Copyright declaration
--	Copyright 2012 林博仁(Henry Lin, pika1021@gmail.com)
--智慧財產授權條款：
--	「設計名稱 | Design name」 is part of 「專案名稱 | Project name」
--	「專案名稱 | Project name」 is free software: you can redistribute it and/or modify it under the terms of the GNU Lesser General Public License as published by the Free Software Foundation, either version 3 of the License, or (at your option) any later version.
--	
--	「專案名稱 | Project name」 is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU Lesser General Public License for more details.
--	
--	You should have received a copy of the GNU Lesser General Public License along with 「專案名稱 | Project name」.  If not, see <http://www.gnu.org/licenses/>.
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity entity_name is
  port (
		: in std_logic;
		: out std_logic
	);
end entity_name;

architecture architecture_name of entity_name is
	--signal : std_logic;
end architecture;
